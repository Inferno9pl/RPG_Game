<?xml version="1.0"?>
<Knight xmlns:xsi="http://www.w3.org/2001/XMLSchema-instance" xmlns:xsd="http://www.w3.org/2001/XMLSchema">
  <Name>Jack</Name>
  <Life>105</Life>
  <MaxLife>568</MaxLife>
  <Level>44</Level>
  <Strenght>111</Strenght>
  <Agility>10</Agility>
  <Eq>
    <Armors>
      <Armors>
        <Armor>
          <Name>Ciężki pancerz łowcy smoków</Name>
          <Value>20000</Value>
          <MeleeProtection>150</MeleeProtection>
          <ArrowProtection>150</ArrowProtection>
          <FireProtection>100</FireProtection>
          <MagicProtection>50</MagicProtection>
        </Armor>
      </Armors>
    </Armors>
    <Weapons>
      <Weapons>
        <Weapon>
          <Name>Gniew Innosa</Name>
          <Value>4000</Value>
          <Type>74</Type>
          <Damage>140</Damage>
          <Requirement>100</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
        <Weapon>
          <Name>Orkowy miecz wojenny</Name>
          <Value>130</Value>
          <Type>68</Type>
          <Damage>100</Damage>
          <Requirement>120</Requirement>
          <Stat>83</Stat>
        </Weapon>
      </Weapons>
    </Weapons>
    <Items>
      <Items>
        <ItemAndQuantity>
          <Item>
            <Name>esencja lecznicza</Name>
            <Value>26</Value>
            <Type>mikstura</Type>
            <Number>50</Number>
          </Item>
          <Quantity>37</Quantity>
        </ItemAndQuantity>
        <ItemAndQuantity>
          <Item>
            <Name>ekstrakt leczniczy</Name>
            <Value>35</Value>
            <Type>mikstura</Type>
            <Number>70</Number>
          </Item>
          <Quantity>39</Quantity>
        </ItemAndQuantity>
        <ItemAndQuantity>
          <Item>
            <Name>eliksir leczniczy</Name>
            <Value>50</Value>
            <Type>mikstura</Type>
            <Number>100</Number>
          </Item>
          <Quantity>46</Quantity>
        </ItemAndQuantity>
        <ItemAndQuantity>
          <Item>
            <Name>gulasz</Name>
            <Value>8</Value>
            <Type>pożywienie</Type>
            <Number>20</Number>
          </Item>
          <Quantity>4</Quantity>
        </ItemAndQuantity>
        <ItemAndQuantity>
          <Item>
            <Name>śledź</Name>
            <Value>15</Value>
            <Type>pożywienie</Type>
            <Number>20</Number>
          </Item>
          <Quantity>10</Quantity>
        </ItemAndQuantity>
        <ItemAndQuantity>
          <Item>
            <Name>serce lodowego golema</Name>
            <Value>300</Value>
            <Type>trofeum</Type>
            <Number>-1</Number>
          </Item>
          <Quantity>21</Quantity>
        </ItemAndQuantity>
        <ItemAndQuantity>
          <Item>
            <Name>skóra warga</Name>
            <Value>25</Value>
            <Type>skóra</Type>
            <Number>-1</Number>
          </Item>
          <Quantity>29</Quantity>
        </ItemAndQuantity>
        <ItemAndQuantity>
          <Item>
            <Name>smażone mięso</Name>
            <Value>6</Value>
            <Type>pożywienie</Type>
            <Number>12</Number>
          </Item>
          <Quantity>13</Quantity>
        </ItemAndQuantity>
        <ItemAndQuantity>
          <Item>
            <Name>szynka</Name>
            <Value>50</Value>
            <Type>pożywienie</Type>
            <Number>20</Number>
          </Item>
          <Quantity>1</Quantity>
        </ItemAndQuantity>
        <ItemAndQuantity>
          <Item>
            <Name>mięso chrząszcza</Name>
            <Value>10</Value>
            <Type>pożywienie</Type>
            <Number>10</Number>
          </Item>
          <Quantity>2</Quantity>
        </ItemAndQuantity>
        <ItemAndQuantity>
          <Item>
            <Name>zupa rybna</Name>
            <Value>20</Value>
            <Type>pożywienie</Type>
            <Number>10</Number>
          </Item>
          <Quantity>1</Quantity>
        </ItemAndQuantity>
        <ItemAndQuantity>
          <Item>
            <Name>barania kiełbasa</Name>
            <Value>9</Value>
            <Type>pożywienie</Type>
            <Number>12</Number>
          </Item>
          <Quantity>6</Quantity>
        </ItemAndQuantity>
      </Items>
    </Items>
    <Gold>165402</Gold>
    <EquippedArmorIndex>0</EquippedArmorIndex>
    <EquippedWeaponIndex>0</EquippedWeaponIndex>
  </Eq>
  <Exp>500010</Exp>
  <SkillPoints>0</SkillPoints>
  <Skill>
    <OneHanded>100</OneHanded>
    <TwoHanded>10</TwoHanded>
    <Bow>10</Bow>
    <Crossbow>10</Crossbow>
  </Skill>
</Knight>