<?xml version="1.0"?>
<Knight xmlns:xsi="http://www.w3.org/2001/XMLSchema-instance" xmlns:xsd="http://www.w3.org/2001/XMLSchema">
  <Name>Wojciech</Name>
  <Life>175</Life>
  <MaxLife>184</MaxLife>
  <Level>12</Level>
  <Strenght>40</Strenght>
  <Agility>10</Agility>
  <Eq>
    <Armors>
      <Armors>
        <Armor>
          <Name>Pancerz Cor Angara</Name>
          <Value>10000</Value>
          <MeleeProtection>100</MeleeProtection>
          <ArrowProtection>100</ArrowProtection>
          <FireProtection>50</FireProtection>
          <MagicProtection>25</MagicProtection>
        </Armor>
      </Armors>
    </Armors>
    <Weapons>
      <Weapons>
        <Weapon>
          <Name>Święty młot</Name>
          <Value>1000</Value>
          <Type>68</Type>
          <Damage>60</Damage>
          <Requirement>10</Requirement>
          <Stat>83</Stat>
        </Weapon>
      </Weapons>
    </Weapons>
    <Items>
      <Items>
        <ItemAndQuantity>
          <Item>
            <Name>smażone mięso</Name>
            <Value>6</Value>
            <Type>pożywienie</Type>
            <Number>12</Number>
          </Item>
          <Quantity>406</Quantity>
        </ItemAndQuantity>
        <ItemAndQuantity>
          <Item>
            <Name>gulasz</Name>
            <Value>8</Value>
            <Type>pożywienie</Type>
            <Number>20</Number>
          </Item>
          <Quantity>133</Quantity>
        </ItemAndQuantity>
        <ItemAndQuantity>
          <Item>
            <Name>żuwaczki pełzacza</Name>
            <Value>15</Value>
            <Type>trofeum</Type>
            <Number>-1</Number>
          </Item>
          <Quantity>3</Quantity>
        </ItemAndQuantity>
        <ItemAndQuantity>
          <Item>
            <Name>płytka pancerza pełzacza</Name>
            <Value>50</Value>
            <Type>trofeum</Type>
            <Number>-1</Number>
          </Item>
          <Quantity>3</Quantity>
        </ItemAndQuantity>
        <ItemAndQuantity>
          <Item>
            <Name>skóra dzika</Name>
            <Value>15</Value>
            <Type>skóra</Type>
            <Number>-1</Number>
          </Item>
          <Quantity>13</Quantity>
        </ItemAndQuantity>
        <ItemAndQuantity>
          <Item>
            <Name>pazury</Name>
            <Value>15</Value>
            <Type>trofeum</Type>
            <Number>-1</Number>
          </Item>
          <Quantity>12</Quantity>
        </ItemAndQuantity>
        <ItemAndQuantity>
          <Item>
            <Name>kieł</Name>
            <Value>15</Value>
            <Type>trofeum</Type>
            <Number>-1</Number>
          </Item>
          <Quantity>8</Quantity>
        </ItemAndQuantity>
        <ItemAndQuantity>
          <Item>
            <Name>skóra topielca</Name>
            <Value>25</Value>
            <Type>skóra</Type>
            <Number>-1</Number>
          </Item>
          <Quantity>4</Quantity>
        </ItemAndQuantity>
        <ItemAndQuantity>
          <Item>
            <Name>szpony topielca</Name>
            <Value>15</Value>
            <Type>trofeum</Type>
            <Number>-1</Number>
          </Item>
          <Quantity>4</Quantity>
        </ItemAndQuantity>
      </Items>
    </Items>
    <Gold>2784</Gold>
    <EquippedArmorIndex>0</EquippedArmorIndex>
    <EquippedWeaponIndex>0</EquippedWeaponIndex>
  </Eq>
  <Exp>39720</Exp>
  <SkillPoints>0</SkillPoints>
  <Skill>
    <OneHanded>10</OneHanded>
    <TwoHanded>64</TwoHanded>
    <Bow>10</Bow>
    <Crossbow>10</Crossbow>
  </Skill>
</Knight>